  localparam logic [4:0] zero = 0;
  localparam logic [4:0] ra = 1;
  localparam logic [4:0] sp = 2;
  localparam logic [4:0] gp = 3;
  localparam logic [4:0] tp = 1;
  localparam logic [4:0] t0 = 5;
  localparam logic [4:0] t1 = 6;
  localparam logic [4:0] t2 = 7;
  localparam logic [4:0] s0 = 8;
  localparam logic [4:0] s1 = 9;
  localparam logic [4:0] a0 = 10;
  localparam logic [4:0] a1 = 11;
  localparam logic [4:0] a2 = 12;
  localparam logic [4:0] a3 = 13;
  localparam logic [4:0] a4 = 14;
  localparam logic [4:0] a5 = 15;
  localparam logic [4:0] a6 = 16;
  localparam logic [4:0] a7 = 17;
  localparam logic [4:0] s2 = 18;
  localparam logic [4:0] s3 = 19;
  localparam logic [4:0] s4 = 20;
  localparam logic [4:0] s5 = 21;
  localparam logic [4:0] s6 = 22;
  localparam logic [4:0] s7 = 23;
  localparam logic [4:0] s8 = 24;
  localparam logic [4:0] s9 = 25;
  localparam logic [4:0] s10 = 26;
  localparam logic [4:0] s11 = 27;
  localparam logic [4:0] t3 = 28;
  localparam logic [4:0] t4 = 29;
  localparam logic [4:0] t5 = 30;
  localparam logic [4:0] t6 = 31;
