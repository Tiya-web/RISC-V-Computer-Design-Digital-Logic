`define E(m) $sformatf("ERROR: %s:%0d: %s", `__FILE__, `__LINE__, m)
